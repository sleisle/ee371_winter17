// nios_system_checkersv3.v

// Generated using ACDS version 14.0 200 at 2017.03.07.23:37:26

`timescale 1 ps / 1 ps
module nios_system_checkersv3 (
		input  wire        clk_clk,             //          clk.clk
		input  wire        reset_reset_n,       //        reset.reset_n
		output wire [7:0]  sendstate_export,    //    sendstate.export
		input  wire [7:0]  receivestate_export, // receivestate.export
		input  wire [7:0]  newdata_export,      //      newdata.export
		input  wire [31:0] row8_in_port,        //         row8.in_port
		output wire [31:0] row8_out_port,       //             .out_port
		input  wire [31:0] row7_in_port,        //         row7.in_port
		output wire [31:0] row7_out_port,       //             .out_port
		input  wire [31:0] row6_in_port,        //         row6.in_port
		output wire [31:0] row6_out_port,       //             .out_port
		input  wire [31:0] row5_in_port,        //         row5.in_port
		output wire [31:0] row5_out_port,       //             .out_port
		input  wire [31:0] row4_in_port,        //         row4.in_port
		output wire [31:0] row4_out_port,       //             .out_port
		input  wire [31:0] row3_in_port,        //         row3.in_port
		output wire [31:0] row3_out_port,       //             .out_port
		input  wire [31:0] row2_in_port,        //         row2.in_port
		output wire [31:0] row2_out_port,       //             .out_port
		input  wire [31:0] row1_in_port,        //         row1.in_port
		output wire [31:0] row1_out_port        //             .out_port
	);

	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [18:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [18:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire  [31:0] mm_interconnect_0_sendstate_s1_writedata;                     // mm_interconnect_0:sendState_s1_writedata -> sendState:writedata
	wire   [1:0] mm_interconnect_0_sendstate_s1_address;                       // mm_interconnect_0:sendState_s1_address -> sendState:address
	wire         mm_interconnect_0_sendstate_s1_chipselect;                    // mm_interconnect_0:sendState_s1_chipselect -> sendState:chipselect
	wire         mm_interconnect_0_sendstate_s1_write;                         // mm_interconnect_0:sendState_s1_write -> sendState:write_n
	wire  [31:0] mm_interconnect_0_sendstate_s1_readdata;                      // sendState:readdata -> mm_interconnect_0:sendState_s1_readdata
	wire   [1:0] mm_interconnect_0_receivestate_s1_address;                    // mm_interconnect_0:receiveState_s1_address -> receiveState:address
	wire  [31:0] mm_interconnect_0_receivestate_s1_readdata;                   // receiveState:readdata -> mm_interconnect_0:receiveState_s1_readdata
	wire   [1:0] mm_interconnect_0_newdata_s1_address;                         // mm_interconnect_0:newData_s1_address -> newData:address
	wire  [31:0] mm_interconnect_0_newdata_s1_readdata;                        // newData:readdata -> mm_interconnect_0:newData_s1_readdata
	wire  [31:0] mm_interconnect_0_row8_s1_writedata;                          // mm_interconnect_0:row8_s1_writedata -> row8:writedata
	wire   [2:0] mm_interconnect_0_row8_s1_address;                            // mm_interconnect_0:row8_s1_address -> row8:address
	wire         mm_interconnect_0_row8_s1_chipselect;                         // mm_interconnect_0:row8_s1_chipselect -> row8:chipselect
	wire         mm_interconnect_0_row8_s1_write;                              // mm_interconnect_0:row8_s1_write -> row8:write_n
	wire  [31:0] mm_interconnect_0_row8_s1_readdata;                           // row8:readdata -> mm_interconnect_0:row8_s1_readdata
	wire  [31:0] mm_interconnect_0_row7_s1_writedata;                          // mm_interconnect_0:row7_s1_writedata -> row7:writedata
	wire   [2:0] mm_interconnect_0_row7_s1_address;                            // mm_interconnect_0:row7_s1_address -> row7:address
	wire         mm_interconnect_0_row7_s1_chipselect;                         // mm_interconnect_0:row7_s1_chipselect -> row7:chipselect
	wire         mm_interconnect_0_row7_s1_write;                              // mm_interconnect_0:row7_s1_write -> row7:write_n
	wire  [31:0] mm_interconnect_0_row7_s1_readdata;                           // row7:readdata -> mm_interconnect_0:row7_s1_readdata
	wire  [31:0] mm_interconnect_0_row6_s1_writedata;                          // mm_interconnect_0:row6_s1_writedata -> row6:writedata
	wire   [2:0] mm_interconnect_0_row6_s1_address;                            // mm_interconnect_0:row6_s1_address -> row6:address
	wire         mm_interconnect_0_row6_s1_chipselect;                         // mm_interconnect_0:row6_s1_chipselect -> row6:chipselect
	wire         mm_interconnect_0_row6_s1_write;                              // mm_interconnect_0:row6_s1_write -> row6:write_n
	wire  [31:0] mm_interconnect_0_row6_s1_readdata;                           // row6:readdata -> mm_interconnect_0:row6_s1_readdata
	wire  [31:0] mm_interconnect_0_row5_s1_writedata;                          // mm_interconnect_0:row5_s1_writedata -> row5:writedata
	wire   [2:0] mm_interconnect_0_row5_s1_address;                            // mm_interconnect_0:row5_s1_address -> row5:address
	wire         mm_interconnect_0_row5_s1_chipselect;                         // mm_interconnect_0:row5_s1_chipselect -> row5:chipselect
	wire         mm_interconnect_0_row5_s1_write;                              // mm_interconnect_0:row5_s1_write -> row5:write_n
	wire  [31:0] mm_interconnect_0_row5_s1_readdata;                           // row5:readdata -> mm_interconnect_0:row5_s1_readdata
	wire  [31:0] mm_interconnect_0_row4_s1_writedata;                          // mm_interconnect_0:row4_s1_writedata -> row4:writedata
	wire   [2:0] mm_interconnect_0_row4_s1_address;                            // mm_interconnect_0:row4_s1_address -> row4:address
	wire         mm_interconnect_0_row4_s1_chipselect;                         // mm_interconnect_0:row4_s1_chipselect -> row4:chipselect
	wire         mm_interconnect_0_row4_s1_write;                              // mm_interconnect_0:row4_s1_write -> row4:write_n
	wire  [31:0] mm_interconnect_0_row4_s1_readdata;                           // row4:readdata -> mm_interconnect_0:row4_s1_readdata
	wire  [31:0] mm_interconnect_0_row3_s1_writedata;                          // mm_interconnect_0:row3_s1_writedata -> row3:writedata
	wire   [2:0] mm_interconnect_0_row3_s1_address;                            // mm_interconnect_0:row3_s1_address -> row3:address
	wire         mm_interconnect_0_row3_s1_chipselect;                         // mm_interconnect_0:row3_s1_chipselect -> row3:chipselect
	wire         mm_interconnect_0_row3_s1_write;                              // mm_interconnect_0:row3_s1_write -> row3:write_n
	wire  [31:0] mm_interconnect_0_row3_s1_readdata;                           // row3:readdata -> mm_interconnect_0:row3_s1_readdata
	wire  [31:0] mm_interconnect_0_row2_s1_writedata;                          // mm_interconnect_0:row2_s1_writedata -> row2:writedata
	wire   [2:0] mm_interconnect_0_row2_s1_address;                            // mm_interconnect_0:row2_s1_address -> row2:address
	wire         mm_interconnect_0_row2_s1_chipselect;                         // mm_interconnect_0:row2_s1_chipselect -> row2:chipselect
	wire         mm_interconnect_0_row2_s1_write;                              // mm_interconnect_0:row2_s1_write -> row2:write_n
	wire  [31:0] mm_interconnect_0_row2_s1_readdata;                           // row2:readdata -> mm_interconnect_0:row2_s1_readdata
	wire  [31:0] mm_interconnect_0_row1_s1_writedata;                          // mm_interconnect_0:row1_s1_writedata -> row1:writedata
	wire   [2:0] mm_interconnect_0_row1_s1_address;                            // mm_interconnect_0:row1_s1_address -> row1:address
	wire         mm_interconnect_0_row1_s1_chipselect;                         // mm_interconnect_0:row1_s1_chipselect -> row1:chipselect
	wire         mm_interconnect_0_row1_s1_write;                              // mm_interconnect_0:row1_s1_write -> row1:write_n
	wire  [31:0] mm_interconnect_0_row1_s1_readdata;                           // row1:readdata -> mm_interconnect_0:row1_s1_readdata
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, newData:reset_n, nios2_qsys_0:reset_n, onchip_memory2_0:reset, receiveState:reset_n, row1:reset_n, row2:reset_n, row3:reset_n, row4:reset_n, row5:reset_n, row6:reset_n, row7:reset_n, row8:reset_n, rst_translator:in_reset, sendState:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios_system_checkersv3_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_checkersv3_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	nios_system_checkersv3_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	nios_system_checkersv3_sendState sendstate (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_sendstate_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sendstate_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sendstate_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sendstate_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sendstate_s1_readdata),   //                    .readdata
		.out_port   (sendstate_export)                           // external_connection.export
	);

	nios_system_checkersv3_receiveState receivestate (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_receivestate_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receivestate_s1_readdata), //                    .readdata
		.in_port  (receivestate_export)                         // external_connection.export
	);

	nios_system_checkersv3_receiveState newdata (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_newdata_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_newdata_s1_readdata), //                    .readdata
		.in_port  (newdata_export)                         // external_connection.export
	);

	nios_system_checkersv3_row8 row8 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_row8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row8_s1_readdata),   //                    .readdata
		.in_port    (row8_in_port),                         // external_connection.export
		.out_port   (row8_out_port)                         //                    .export
	);

	nios_system_checkersv3_row8 row7 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_row7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row7_s1_readdata),   //                    .readdata
		.in_port    (row7_in_port),                         // external_connection.export
		.out_port   (row7_out_port)                         //                    .export
	);

	nios_system_checkersv3_row8 row6 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_row6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row6_s1_readdata),   //                    .readdata
		.in_port    (row6_in_port),                         // external_connection.export
		.out_port   (row6_out_port)                         //                    .export
	);

	nios_system_checkersv3_row8 row5 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_row5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row5_s1_readdata),   //                    .readdata
		.in_port    (row5_in_port),                         // external_connection.export
		.out_port   (row5_out_port)                         //                    .export
	);

	nios_system_checkersv3_row8 row4 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_row4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row4_s1_readdata),   //                    .readdata
		.in_port    (row4_in_port),                         // external_connection.export
		.out_port   (row4_out_port)                         //                    .export
	);

	nios_system_checkersv3_row8 row3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_row3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row3_s1_readdata),   //                    .readdata
		.in_port    (row3_in_port),                         // external_connection.export
		.out_port   (row3_out_port)                         //                    .export
	);

	nios_system_checkersv3_row8 row2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_row2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row2_s1_readdata),   //                    .readdata
		.in_port    (row2_in_port),                         // external_connection.export
		.out_port   (row2_out_port)                         //                    .export
	);

	nios_system_checkersv3_row8 row1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_row1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row1_s1_readdata),   //                    .readdata
		.in_port    (row1_in_port),                         // external_connection.export
		.out_port   (row1_out_port)                         //                    .export
	);

	nios_system_checkersv3_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.newData_s1_address                               (mm_interconnect_0_newdata_s1_address),                         //                                 newData_s1.address
		.newData_s1_readdata                              (mm_interconnect_0_newdata_s1_readdata),                        //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                           .clken
		.receiveState_s1_address                          (mm_interconnect_0_receivestate_s1_address),                    //                            receiveState_s1.address
		.receiveState_s1_readdata                         (mm_interconnect_0_receivestate_s1_readdata),                   //                                           .readdata
		.row1_s1_address                                  (mm_interconnect_0_row1_s1_address),                            //                                    row1_s1.address
		.row1_s1_write                                    (mm_interconnect_0_row1_s1_write),                              //                                           .write
		.row1_s1_readdata                                 (mm_interconnect_0_row1_s1_readdata),                           //                                           .readdata
		.row1_s1_writedata                                (mm_interconnect_0_row1_s1_writedata),                          //                                           .writedata
		.row1_s1_chipselect                               (mm_interconnect_0_row1_s1_chipselect),                         //                                           .chipselect
		.row2_s1_address                                  (mm_interconnect_0_row2_s1_address),                            //                                    row2_s1.address
		.row2_s1_write                                    (mm_interconnect_0_row2_s1_write),                              //                                           .write
		.row2_s1_readdata                                 (mm_interconnect_0_row2_s1_readdata),                           //                                           .readdata
		.row2_s1_writedata                                (mm_interconnect_0_row2_s1_writedata),                          //                                           .writedata
		.row2_s1_chipselect                               (mm_interconnect_0_row2_s1_chipselect),                         //                                           .chipselect
		.row3_s1_address                                  (mm_interconnect_0_row3_s1_address),                            //                                    row3_s1.address
		.row3_s1_write                                    (mm_interconnect_0_row3_s1_write),                              //                                           .write
		.row3_s1_readdata                                 (mm_interconnect_0_row3_s1_readdata),                           //                                           .readdata
		.row3_s1_writedata                                (mm_interconnect_0_row3_s1_writedata),                          //                                           .writedata
		.row3_s1_chipselect                               (mm_interconnect_0_row3_s1_chipselect),                         //                                           .chipselect
		.row4_s1_address                                  (mm_interconnect_0_row4_s1_address),                            //                                    row4_s1.address
		.row4_s1_write                                    (mm_interconnect_0_row4_s1_write),                              //                                           .write
		.row4_s1_readdata                                 (mm_interconnect_0_row4_s1_readdata),                           //                                           .readdata
		.row4_s1_writedata                                (mm_interconnect_0_row4_s1_writedata),                          //                                           .writedata
		.row4_s1_chipselect                               (mm_interconnect_0_row4_s1_chipselect),                         //                                           .chipselect
		.row5_s1_address                                  (mm_interconnect_0_row5_s1_address),                            //                                    row5_s1.address
		.row5_s1_write                                    (mm_interconnect_0_row5_s1_write),                              //                                           .write
		.row5_s1_readdata                                 (mm_interconnect_0_row5_s1_readdata),                           //                                           .readdata
		.row5_s1_writedata                                (mm_interconnect_0_row5_s1_writedata),                          //                                           .writedata
		.row5_s1_chipselect                               (mm_interconnect_0_row5_s1_chipselect),                         //                                           .chipselect
		.row6_s1_address                                  (mm_interconnect_0_row6_s1_address),                            //                                    row6_s1.address
		.row6_s1_write                                    (mm_interconnect_0_row6_s1_write),                              //                                           .write
		.row6_s1_readdata                                 (mm_interconnect_0_row6_s1_readdata),                           //                                           .readdata
		.row6_s1_writedata                                (mm_interconnect_0_row6_s1_writedata),                          //                                           .writedata
		.row6_s1_chipselect                               (mm_interconnect_0_row6_s1_chipselect),                         //                                           .chipselect
		.row7_s1_address                                  (mm_interconnect_0_row7_s1_address),                            //                                    row7_s1.address
		.row7_s1_write                                    (mm_interconnect_0_row7_s1_write),                              //                                           .write
		.row7_s1_readdata                                 (mm_interconnect_0_row7_s1_readdata),                           //                                           .readdata
		.row7_s1_writedata                                (mm_interconnect_0_row7_s1_writedata),                          //                                           .writedata
		.row7_s1_chipselect                               (mm_interconnect_0_row7_s1_chipselect),                         //                                           .chipselect
		.row8_s1_address                                  (mm_interconnect_0_row8_s1_address),                            //                                    row8_s1.address
		.row8_s1_write                                    (mm_interconnect_0_row8_s1_write),                              //                                           .write
		.row8_s1_readdata                                 (mm_interconnect_0_row8_s1_readdata),                           //                                           .readdata
		.row8_s1_writedata                                (mm_interconnect_0_row8_s1_writedata),                          //                                           .writedata
		.row8_s1_chipselect                               (mm_interconnect_0_row8_s1_chipselect),                         //                                           .chipselect
		.sendState_s1_address                             (mm_interconnect_0_sendstate_s1_address),                       //                               sendState_s1.address
		.sendState_s1_write                               (mm_interconnect_0_sendstate_s1_write),                         //                                           .write
		.sendState_s1_readdata                            (mm_interconnect_0_sendstate_s1_readdata),                      //                                           .readdata
		.sendState_s1_writedata                           (mm_interconnect_0_sendstate_s1_writedata),                     //                                           .writedata
		.sendState_s1_chipselect                          (mm_interconnect_0_sendstate_s1_chipselect)                     //                                           .chipselect
	);

	nios_system_checkersv3_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
