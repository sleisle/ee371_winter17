// nios_system_checkersv4.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module nios_system_checkersv4 (
		input  wire        clk_clk,             //          clk.clk
		input  wire [7:0]  newdata_export,      //      newdata.export
		input  wire [7:0]  receivestate_export, // receivestate.export
		input  wire        reset_reset_n,       //        reset.reset_n
		input  wire [31:0] row1in_export,       //       row1in.export
		output wire [31:0] row1out_export,      //      row1out.export
		input  wire [31:0] row2in_export,       //       row2in.export
		output wire [31:0] row2out_export,      //      row2out.export
		input  wire [31:0] row3in_export,       //       row3in.export
		output wire [31:0] row3out_export,      //      row3out.export
		input  wire [31:0] row4in_export,       //       row4in.export
		output wire [31:0] row4out_export,      //      row4out.export
		input  wire [31:0] row5in_export,       //       row5in.export
		output wire [31:0] row5out_export,      //      row5out.export
		input  wire [31:0] row6in_export,       //       row6in.export
		output wire [31:0] row6out_export,      //      row6out.export
		input  wire [31:0] row7in_export,       //       row7in.export
		output wire [31:0] row7out_export,      //      row7out.export
		input  wire [31:0] row8in_export,       //       row8in.export
		output wire [31:0] row8out_export,      //      row8out.export
		output wire [7:0]  sendstate_export     //    sendstate.export
	);

	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [18:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [18:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sendstate_s1_chipselect;                    // mm_interconnect_0:sendState_s1_chipselect -> sendState:chipselect
	wire  [31:0] mm_interconnect_0_sendstate_s1_readdata;                      // sendState:readdata -> mm_interconnect_0:sendState_s1_readdata
	wire   [1:0] mm_interconnect_0_sendstate_s1_address;                       // mm_interconnect_0:sendState_s1_address -> sendState:address
	wire         mm_interconnect_0_sendstate_s1_write;                         // mm_interconnect_0:sendState_s1_write -> sendState:write_n
	wire  [31:0] mm_interconnect_0_sendstate_s1_writedata;                     // mm_interconnect_0:sendState_s1_writedata -> sendState:writedata
	wire  [31:0] mm_interconnect_0_receivestate_s1_readdata;                   // receiveState:readdata -> mm_interconnect_0:receiveState_s1_readdata
	wire   [1:0] mm_interconnect_0_receivestate_s1_address;                    // mm_interconnect_0:receiveState_s1_address -> receiveState:address
	wire  [31:0] mm_interconnect_0_newdata_s1_readdata;                        // newData:readdata -> mm_interconnect_0:newData_s1_readdata
	wire   [1:0] mm_interconnect_0_newdata_s1_address;                         // mm_interconnect_0:newData_s1_address -> newData:address
	wire         mm_interconnect_0_row8out_s1_chipselect;                      // mm_interconnect_0:row8out_s1_chipselect -> row8out:chipselect
	wire  [31:0] mm_interconnect_0_row8out_s1_readdata;                        // row8out:readdata -> mm_interconnect_0:row8out_s1_readdata
	wire   [2:0] mm_interconnect_0_row8out_s1_address;                         // mm_interconnect_0:row8out_s1_address -> row8out:address
	wire         mm_interconnect_0_row8out_s1_write;                           // mm_interconnect_0:row8out_s1_write -> row8out:write_n
	wire  [31:0] mm_interconnect_0_row8out_s1_writedata;                       // mm_interconnect_0:row8out_s1_writedata -> row8out:writedata
	wire         mm_interconnect_0_row7out_s1_chipselect;                      // mm_interconnect_0:row7out_s1_chipselect -> row7out:chipselect
	wire  [31:0] mm_interconnect_0_row7out_s1_readdata;                        // row7out:readdata -> mm_interconnect_0:row7out_s1_readdata
	wire   [2:0] mm_interconnect_0_row7out_s1_address;                         // mm_interconnect_0:row7out_s1_address -> row7out:address
	wire         mm_interconnect_0_row7out_s1_write;                           // mm_interconnect_0:row7out_s1_write -> row7out:write_n
	wire  [31:0] mm_interconnect_0_row7out_s1_writedata;                       // mm_interconnect_0:row7out_s1_writedata -> row7out:writedata
	wire         mm_interconnect_0_row6out_s1_chipselect;                      // mm_interconnect_0:row6out_s1_chipselect -> row6out:chipselect
	wire  [31:0] mm_interconnect_0_row6out_s1_readdata;                        // row6out:readdata -> mm_interconnect_0:row6out_s1_readdata
	wire   [2:0] mm_interconnect_0_row6out_s1_address;                         // mm_interconnect_0:row6out_s1_address -> row6out:address
	wire         mm_interconnect_0_row6out_s1_write;                           // mm_interconnect_0:row6out_s1_write -> row6out:write_n
	wire  [31:0] mm_interconnect_0_row6out_s1_writedata;                       // mm_interconnect_0:row6out_s1_writedata -> row6out:writedata
	wire         mm_interconnect_0_row5out_s1_chipselect;                      // mm_interconnect_0:row5out_s1_chipselect -> row5out:chipselect
	wire  [31:0] mm_interconnect_0_row5out_s1_readdata;                        // row5out:readdata -> mm_interconnect_0:row5out_s1_readdata
	wire   [2:0] mm_interconnect_0_row5out_s1_address;                         // mm_interconnect_0:row5out_s1_address -> row5out:address
	wire         mm_interconnect_0_row5out_s1_write;                           // mm_interconnect_0:row5out_s1_write -> row5out:write_n
	wire  [31:0] mm_interconnect_0_row5out_s1_writedata;                       // mm_interconnect_0:row5out_s1_writedata -> row5out:writedata
	wire         mm_interconnect_0_row4out_s1_chipselect;                      // mm_interconnect_0:row4out_s1_chipselect -> row4out:chipselect
	wire  [31:0] mm_interconnect_0_row4out_s1_readdata;                        // row4out:readdata -> mm_interconnect_0:row4out_s1_readdata
	wire   [2:0] mm_interconnect_0_row4out_s1_address;                         // mm_interconnect_0:row4out_s1_address -> row4out:address
	wire         mm_interconnect_0_row4out_s1_write;                           // mm_interconnect_0:row4out_s1_write -> row4out:write_n
	wire  [31:0] mm_interconnect_0_row4out_s1_writedata;                       // mm_interconnect_0:row4out_s1_writedata -> row4out:writedata
	wire         mm_interconnect_0_row3out_s1_chipselect;                      // mm_interconnect_0:row3out_s1_chipselect -> row3out:chipselect
	wire  [31:0] mm_interconnect_0_row3out_s1_readdata;                        // row3out:readdata -> mm_interconnect_0:row3out_s1_readdata
	wire   [2:0] mm_interconnect_0_row3out_s1_address;                         // mm_interconnect_0:row3out_s1_address -> row3out:address
	wire         mm_interconnect_0_row3out_s1_write;                           // mm_interconnect_0:row3out_s1_write -> row3out:write_n
	wire  [31:0] mm_interconnect_0_row3out_s1_writedata;                       // mm_interconnect_0:row3out_s1_writedata -> row3out:writedata
	wire         mm_interconnect_0_row2out_s1_chipselect;                      // mm_interconnect_0:row2out_s1_chipselect -> row2out:chipselect
	wire  [31:0] mm_interconnect_0_row2out_s1_readdata;                        // row2out:readdata -> mm_interconnect_0:row2out_s1_readdata
	wire   [2:0] mm_interconnect_0_row2out_s1_address;                         // mm_interconnect_0:row2out_s1_address -> row2out:address
	wire         mm_interconnect_0_row2out_s1_write;                           // mm_interconnect_0:row2out_s1_write -> row2out:write_n
	wire  [31:0] mm_interconnect_0_row2out_s1_writedata;                       // mm_interconnect_0:row2out_s1_writedata -> row2out:writedata
	wire         mm_interconnect_0_row1out_s1_chipselect;                      // mm_interconnect_0:row1out_s1_chipselect -> row1out:chipselect
	wire  [31:0] mm_interconnect_0_row1out_s1_readdata;                        // row1out:readdata -> mm_interconnect_0:row1out_s1_readdata
	wire   [2:0] mm_interconnect_0_row1out_s1_address;                         // mm_interconnect_0:row1out_s1_address -> row1out:address
	wire         mm_interconnect_0_row1out_s1_write;                           // mm_interconnect_0:row1out_s1_write -> row1out:write_n
	wire  [31:0] mm_interconnect_0_row1out_s1_writedata;                       // mm_interconnect_0:row1out_s1_writedata -> row1out:writedata
	wire  [31:0] mm_interconnect_0_row8in_s1_readdata;                         // row8in:readdata -> mm_interconnect_0:row8in_s1_readdata
	wire   [1:0] mm_interconnect_0_row8in_s1_address;                          // mm_interconnect_0:row8in_s1_address -> row8in:address
	wire  [31:0] mm_interconnect_0_row7in_s1_readdata;                         // row7in:readdata -> mm_interconnect_0:row7in_s1_readdata
	wire   [1:0] mm_interconnect_0_row7in_s1_address;                          // mm_interconnect_0:row7in_s1_address -> row7in:address
	wire  [31:0] mm_interconnect_0_row6in_s1_readdata;                         // row6in:readdata -> mm_interconnect_0:row6in_s1_readdata
	wire   [1:0] mm_interconnect_0_row6in_s1_address;                          // mm_interconnect_0:row6in_s1_address -> row6in:address
	wire  [31:0] mm_interconnect_0_row5in_s1_readdata;                         // row5in:readdata -> mm_interconnect_0:row5in_s1_readdata
	wire   [1:0] mm_interconnect_0_row5in_s1_address;                          // mm_interconnect_0:row5in_s1_address -> row5in:address
	wire  [31:0] mm_interconnect_0_row4in_s1_readdata;                         // row4in:readdata -> mm_interconnect_0:row4in_s1_readdata
	wire   [1:0] mm_interconnect_0_row4in_s1_address;                          // mm_interconnect_0:row4in_s1_address -> row4in:address
	wire  [31:0] mm_interconnect_0_row3in_s1_readdata;                         // row3in:readdata -> mm_interconnect_0:row3in_s1_readdata
	wire   [1:0] mm_interconnect_0_row3in_s1_address;                          // mm_interconnect_0:row3in_s1_address -> row3in:address
	wire  [31:0] mm_interconnect_0_row2in_s1_readdata;                         // row2in:readdata -> mm_interconnect_0:row2in_s1_readdata
	wire   [1:0] mm_interconnect_0_row2in_s1_address;                          // mm_interconnect_0:row2in_s1_address -> row2in:address
	wire  [31:0] mm_interconnect_0_row1in_s1_readdata;                         // row1in:readdata -> mm_interconnect_0:row1in_s1_readdata
	wire   [1:0] mm_interconnect_0_row1in_s1_address;                          // mm_interconnect_0:row1in_s1_address -> row1in:address
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, newData:reset_n, nios2_qsys_0:reset_n, onchip_memory2_0:reset, receiveState:reset_n, row1in:reset_n, row1out:reset_n, row2in:reset_n, row2out:reset_n, row3in:reset_n, row3out:reset_n, row4in:reset_n, row4out:reset_n, row5in:reset_n, row5out:reset_n, row6in:reset_n, row6out:reset_n, row7in:reset_n, row7out:reset_n, row8in:reset_n, row8out:reset_n, rst_translator:in_reset, sendState:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios_system_checkersv4_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_checkersv4_newData newdata (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_newdata_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_newdata_s1_readdata), //                    .readdata
		.in_port  (newdata_export)                         // external_connection.export
	);

	nios_system_checkersv4_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	nios_system_checkersv4_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	nios_system_checkersv4_newData receivestate (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_receivestate_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receivestate_s1_readdata), //                    .readdata
		.in_port  (receivestate_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1in row1in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_row1in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_row1in_s1_readdata), //                    .readdata
		.in_port  (row1in_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1out row1out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_row1out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row1out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row1out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row1out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row1out_s1_readdata),   //                    .readdata
		.out_port   (row1out_export)                           // external_connection.export
	);

	nios_system_checkersv4_row1in row2in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_row2in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_row2in_s1_readdata), //                    .readdata
		.in_port  (row2in_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1out row2out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_row2out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row2out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row2out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row2out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row2out_s1_readdata),   //                    .readdata
		.out_port   (row2out_export)                           // external_connection.export
	);

	nios_system_checkersv4_row1in row3in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_row3in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_row3in_s1_readdata), //                    .readdata
		.in_port  (row3in_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1out row3out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_row3out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row3out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row3out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row3out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row3out_s1_readdata),   //                    .readdata
		.out_port   (row3out_export)                           // external_connection.export
	);

	nios_system_checkersv4_row1in row4in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_row4in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_row4in_s1_readdata), //                    .readdata
		.in_port  (row4in_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1out row4out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_row4out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row4out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row4out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row4out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row4out_s1_readdata),   //                    .readdata
		.out_port   (row4out_export)                           // external_connection.export
	);

	nios_system_checkersv4_row1in row5in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_row5in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_row5in_s1_readdata), //                    .readdata
		.in_port  (row5in_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1out row5out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_row5out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row5out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row5out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row5out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row5out_s1_readdata),   //                    .readdata
		.out_port   (row5out_export)                           // external_connection.export
	);

	nios_system_checkersv4_row1in row6in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_row6in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_row6in_s1_readdata), //                    .readdata
		.in_port  (row6in_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1out row6out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_row6out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row6out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row6out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row6out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row6out_s1_readdata),   //                    .readdata
		.out_port   (row6out_export)                           // external_connection.export
	);

	nios_system_checkersv4_row1in row7in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_row7in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_row7in_s1_readdata), //                    .readdata
		.in_port  (row7in_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1out row7out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_row7out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row7out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row7out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row7out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row7out_s1_readdata),   //                    .readdata
		.out_port   (row7out_export)                           // external_connection.export
	);

	nios_system_checkersv4_row1in row8in (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_row8in_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_row8in_s1_readdata), //                    .readdata
		.in_port  (row8in_export)                         // external_connection.export
	);

	nios_system_checkersv4_row1out row8out (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_row8out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_row8out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_row8out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_row8out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_row8out_s1_readdata),   //                    .readdata
		.out_port   (row8out_export)                           // external_connection.export
	);

	nios_system_checkersv4_sendState sendstate (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_sendstate_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sendstate_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sendstate_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sendstate_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sendstate_s1_readdata),   //                    .readdata
		.out_port   (sendstate_export)                           // external_connection.export
	);

	nios_system_checkersv4_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                    (clk_clk),                                                      //                                  clk_0_clk.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                 (nios2_qsys_0_data_master_address),                             //                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest             (nios2_qsys_0_data_master_waitrequest),                         //                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable              (nios2_qsys_0_data_master_byteenable),                          //                                           .byteenable
		.nios2_qsys_0_data_master_read                    (nios2_qsys_0_data_master_read),                                //                                           .read
		.nios2_qsys_0_data_master_readdata                (nios2_qsys_0_data_master_readdata),                            //                                           .readdata
		.nios2_qsys_0_data_master_write                   (nios2_qsys_0_data_master_write),                               //                                           .write
		.nios2_qsys_0_data_master_writedata               (nios2_qsys_0_data_master_writedata),                           //                                           .writedata
		.nios2_qsys_0_data_master_debugaccess             (nios2_qsys_0_data_master_debugaccess),                         //                                           .debugaccess
		.nios2_qsys_0_instruction_master_address          (nios2_qsys_0_instruction_master_address),                      //            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest      (nios2_qsys_0_instruction_master_waitrequest),                  //                                           .waitrequest
		.nios2_qsys_0_instruction_master_read             (nios2_qsys_0_instruction_master_read),                         //                                           .read
		.nios2_qsys_0_instruction_master_readdata         (nios2_qsys_0_instruction_master_readdata),                     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_address            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //              jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                           .write
		.jtag_uart_0_avalon_jtag_slave_read               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                           .read
		.jtag_uart_0_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                           .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                           .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                           .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                           .chipselect
		.newData_s1_address                               (mm_interconnect_0_newdata_s1_address),                         //                                 newData_s1.address
		.newData_s1_readdata                              (mm_interconnect_0_newdata_s1_readdata),                        //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_address           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //             nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                           .write
		.nios2_qsys_0_jtag_debug_module_read              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                           .read
		.nios2_qsys_0_jtag_debug_module_readdata          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                           .readdata
		.nios2_qsys_0_jtag_debug_module_writedata         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                           .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                           .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                           .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                           .debugaccess
		.onchip_memory2_0_s1_address                      (mm_interconnect_0_onchip_memory2_0_s1_address),                //                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                        (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                           .write
		.onchip_memory2_0_s1_readdata                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                           .readdata
		.onchip_memory2_0_s1_writedata                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                           .writedata
		.onchip_memory2_0_s1_byteenable                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                           .byteenable
		.onchip_memory2_0_s1_chipselect                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                           .chipselect
		.onchip_memory2_0_s1_clken                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                           .clken
		.receiveState_s1_address                          (mm_interconnect_0_receivestate_s1_address),                    //                            receiveState_s1.address
		.receiveState_s1_readdata                         (mm_interconnect_0_receivestate_s1_readdata),                   //                                           .readdata
		.row1in_s1_address                                (mm_interconnect_0_row1in_s1_address),                          //                                  row1in_s1.address
		.row1in_s1_readdata                               (mm_interconnect_0_row1in_s1_readdata),                         //                                           .readdata
		.row1out_s1_address                               (mm_interconnect_0_row1out_s1_address),                         //                                 row1out_s1.address
		.row1out_s1_write                                 (mm_interconnect_0_row1out_s1_write),                           //                                           .write
		.row1out_s1_readdata                              (mm_interconnect_0_row1out_s1_readdata),                        //                                           .readdata
		.row1out_s1_writedata                             (mm_interconnect_0_row1out_s1_writedata),                       //                                           .writedata
		.row1out_s1_chipselect                            (mm_interconnect_0_row1out_s1_chipselect),                      //                                           .chipselect
		.row2in_s1_address                                (mm_interconnect_0_row2in_s1_address),                          //                                  row2in_s1.address
		.row2in_s1_readdata                               (mm_interconnect_0_row2in_s1_readdata),                         //                                           .readdata
		.row2out_s1_address                               (mm_interconnect_0_row2out_s1_address),                         //                                 row2out_s1.address
		.row2out_s1_write                                 (mm_interconnect_0_row2out_s1_write),                           //                                           .write
		.row2out_s1_readdata                              (mm_interconnect_0_row2out_s1_readdata),                        //                                           .readdata
		.row2out_s1_writedata                             (mm_interconnect_0_row2out_s1_writedata),                       //                                           .writedata
		.row2out_s1_chipselect                            (mm_interconnect_0_row2out_s1_chipselect),                      //                                           .chipselect
		.row3in_s1_address                                (mm_interconnect_0_row3in_s1_address),                          //                                  row3in_s1.address
		.row3in_s1_readdata                               (mm_interconnect_0_row3in_s1_readdata),                         //                                           .readdata
		.row3out_s1_address                               (mm_interconnect_0_row3out_s1_address),                         //                                 row3out_s1.address
		.row3out_s1_write                                 (mm_interconnect_0_row3out_s1_write),                           //                                           .write
		.row3out_s1_readdata                              (mm_interconnect_0_row3out_s1_readdata),                        //                                           .readdata
		.row3out_s1_writedata                             (mm_interconnect_0_row3out_s1_writedata),                       //                                           .writedata
		.row3out_s1_chipselect                            (mm_interconnect_0_row3out_s1_chipselect),                      //                                           .chipselect
		.row4in_s1_address                                (mm_interconnect_0_row4in_s1_address),                          //                                  row4in_s1.address
		.row4in_s1_readdata                               (mm_interconnect_0_row4in_s1_readdata),                         //                                           .readdata
		.row4out_s1_address                               (mm_interconnect_0_row4out_s1_address),                         //                                 row4out_s1.address
		.row4out_s1_write                                 (mm_interconnect_0_row4out_s1_write),                           //                                           .write
		.row4out_s1_readdata                              (mm_interconnect_0_row4out_s1_readdata),                        //                                           .readdata
		.row4out_s1_writedata                             (mm_interconnect_0_row4out_s1_writedata),                       //                                           .writedata
		.row4out_s1_chipselect                            (mm_interconnect_0_row4out_s1_chipselect),                      //                                           .chipselect
		.row5in_s1_address                                (mm_interconnect_0_row5in_s1_address),                          //                                  row5in_s1.address
		.row5in_s1_readdata                               (mm_interconnect_0_row5in_s1_readdata),                         //                                           .readdata
		.row5out_s1_address                               (mm_interconnect_0_row5out_s1_address),                         //                                 row5out_s1.address
		.row5out_s1_write                                 (mm_interconnect_0_row5out_s1_write),                           //                                           .write
		.row5out_s1_readdata                              (mm_interconnect_0_row5out_s1_readdata),                        //                                           .readdata
		.row5out_s1_writedata                             (mm_interconnect_0_row5out_s1_writedata),                       //                                           .writedata
		.row5out_s1_chipselect                            (mm_interconnect_0_row5out_s1_chipselect),                      //                                           .chipselect
		.row6in_s1_address                                (mm_interconnect_0_row6in_s1_address),                          //                                  row6in_s1.address
		.row6in_s1_readdata                               (mm_interconnect_0_row6in_s1_readdata),                         //                                           .readdata
		.row6out_s1_address                               (mm_interconnect_0_row6out_s1_address),                         //                                 row6out_s1.address
		.row6out_s1_write                                 (mm_interconnect_0_row6out_s1_write),                           //                                           .write
		.row6out_s1_readdata                              (mm_interconnect_0_row6out_s1_readdata),                        //                                           .readdata
		.row6out_s1_writedata                             (mm_interconnect_0_row6out_s1_writedata),                       //                                           .writedata
		.row6out_s1_chipselect                            (mm_interconnect_0_row6out_s1_chipselect),                      //                                           .chipselect
		.row7in_s1_address                                (mm_interconnect_0_row7in_s1_address),                          //                                  row7in_s1.address
		.row7in_s1_readdata                               (mm_interconnect_0_row7in_s1_readdata),                         //                                           .readdata
		.row7out_s1_address                               (mm_interconnect_0_row7out_s1_address),                         //                                 row7out_s1.address
		.row7out_s1_write                                 (mm_interconnect_0_row7out_s1_write),                           //                                           .write
		.row7out_s1_readdata                              (mm_interconnect_0_row7out_s1_readdata),                        //                                           .readdata
		.row7out_s1_writedata                             (mm_interconnect_0_row7out_s1_writedata),                       //                                           .writedata
		.row7out_s1_chipselect                            (mm_interconnect_0_row7out_s1_chipselect),                      //                                           .chipselect
		.row8in_s1_address                                (mm_interconnect_0_row8in_s1_address),                          //                                  row8in_s1.address
		.row8in_s1_readdata                               (mm_interconnect_0_row8in_s1_readdata),                         //                                           .readdata
		.row8out_s1_address                               (mm_interconnect_0_row8out_s1_address),                         //                                 row8out_s1.address
		.row8out_s1_write                                 (mm_interconnect_0_row8out_s1_write),                           //                                           .write
		.row8out_s1_readdata                              (mm_interconnect_0_row8out_s1_readdata),                        //                                           .readdata
		.row8out_s1_writedata                             (mm_interconnect_0_row8out_s1_writedata),                       //                                           .writedata
		.row8out_s1_chipselect                            (mm_interconnect_0_row8out_s1_chipselect),                      //                                           .chipselect
		.sendState_s1_address                             (mm_interconnect_0_sendstate_s1_address),                       //                               sendState_s1.address
		.sendState_s1_write                               (mm_interconnect_0_sendstate_s1_write),                         //                                           .write
		.sendState_s1_readdata                            (mm_interconnect_0_sendstate_s1_readdata),                      //                                           .readdata
		.sendState_s1_writedata                           (mm_interconnect_0_sendstate_s1_writedata),                     //                                           .writedata
		.sendState_s1_chipselect                          (mm_interconnect_0_sendstate_s1_chipselect)                     //                                           .chipselect
	);

	nios_system_checkersv4_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
