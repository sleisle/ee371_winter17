module lockSystem ();

endmodule
